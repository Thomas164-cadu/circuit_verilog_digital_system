module BOBC(
    input inicio;
    
);