module BOBC(
    
);