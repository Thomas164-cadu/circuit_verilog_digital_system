module BO (
    input [15:0] A,
    input [15:0] B,
    input [15:0] C,
    input MO,
    input [7:0] X,
    input clk,
    input LX,
    input RSTX,
    input M1,
    input M2,
    input LH,
    input clkH,
    input RSTH,
    input LS,
    input clkS,
    output [15:0] Pronto 
); 
    
endmodule